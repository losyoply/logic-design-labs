module Comparator_4bits (A, B, A_lt_B, A_gt_B, A_eq_B);
// declare input signals
input [4-1:0] A;
input [4-1:0] B;

// declare output signals
output A_lt_B, A_gt_B, A_eq_B;

// here is your design

endmodule




